module CONCAT (a, b, c, concatout);

//concaternar a, b, c
input [4:0] a;
input [4:0] b;
input [15:0] c;
output [25:0] concatout;

endmodule