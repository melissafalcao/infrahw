module SignExtend(concatout, ext25_32);

	input [25:0]  concatout; 
	output reg[31:0]  ext25_32;

endmodule
