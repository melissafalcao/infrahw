module DeslocamentoBox(Shifter, MUX9out, MUX10out, Shiftout);

	input [1:0] Shifter;
	input [31:0] MUX9out, MUX10out; 
	output [31:0] Shiftout; 

endmodule
