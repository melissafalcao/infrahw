module MUX4(ULAa, pc, mdr, a, MUX4out);

	input [1:0] ULAa; 
	input [31:0] pc, mdr, a; 
	output [31:0] MUX4out;

endmodule
