module GetEndOfB(B, endB);

	input [31:0] B; 
	output [4:0]  endB; 

endmodule
