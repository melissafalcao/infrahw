module MUX5(ULAb, B, ext16_32, reg4, reg1, ext16_32_left_shifted, MUX5out);

	input [2:0] ULAb; 
	input [31:0]  B, ext16_32, reg4, reg1, ext16_32_left_shifted; 
	output [31:0] MUX5out;

endmodule
