module ShiftLeft2(ext16_32, ext16_32_left_shift);

	input [31:0]  ext16_32; 
	output [31:0]  ext16_32_left_shift; 

endmodule
