module MUX1 (MemoryAdress, ext35_32, PC, ulaResult, ext16_32, ULAout, reg253, reg254, reg255, MUX1outMUX1out);

input [2:0]MemoryAdress;
input [31:0] ext35_32, PC, ulaResult, ext16_32, ULAout, reg253, reg254, reg255;
output [31:0] MUX1out;

endmodule

