module UnitExtend(LT, LT32);

	input LT; 
	output [31:0]  LT32; 

endmodule
