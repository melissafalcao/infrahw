module HIeLO(HILOWrite, hi, lo, hiout, loout);

	input HILOWrite;
	input [31:0] hi, lo;  
	output [31:0] hiout, loout; 

endmodule
