module MUX14(mux14, ULAresult, LSout, mux14out);

	input mux14; 
	input [31:0]  ULAresult, LSout; 
	output [31:0]  mux14out;

endmodule
