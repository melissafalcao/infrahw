module CONCAT (rs, rt, immediato, concatout);

//concaternar a, b, c
  input [4:0] rs;
  input [4:0] rt;
  input [15:0] immediato;
output [25:0] concatout;

endmodule
