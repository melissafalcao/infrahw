module pc(PCwrite, mux6OUT, pc) 

input PCwrite;
input [31:0] mux6OUT;
output [31:0] pc;
