module GetShamt(imediato, shamt);

	input [15:0] imediato; 
	output [4:0] shamt;

endmodule
