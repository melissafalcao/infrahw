module MUX14(muux14, ULAresult, LSout, mux14out);

	input muux14; 
	input [31:0]  ULAresult, LSout; 
	output [31:0]  mux14out;

endmodule
