module DIVeMULTI(MDcontrol, a, b, hi, lo);

	input MDcontrol;
	input [31:0] a, b;  //fazer div e multi aqui jogando a saida no hi e lo
	output [31:0] hi, lo; 

endmodule
