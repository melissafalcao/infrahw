module SighLeft2Concat(concatout, pc, SLAC);

	input [25:0] concatout; 
	input [31:0]  pc; 
	output [31:0]  SLAC;

endmodule
