module MUX2 (WriteData, ULAout, LSout, HIout, LOout, Shiftout, LT32, MUX2out)

input [2:0] WriteData;
input [31:0]  ULAout, LSout, HIout, LOout, Shiftout, LT32;
output [31:0] MUX2out;


