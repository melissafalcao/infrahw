module MUX6(PCmux, a, ULAout, SLAC, EPCout, MDRout, ULAresult, MUX6out);

	input [2:0]  PCmux; 
	input [31:0]  a, ULAout, SLAC, EPCout, MDRout, ULAresult; 
	output [31:0]  MUX6out;

endmodule
