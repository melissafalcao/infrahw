module EPC(EPCcontrol, mux4out, EPCout);

	input EPCcontrol; 
	input [31:0]  mux4out; 
	output [31:0] EPCout;

endmodule
