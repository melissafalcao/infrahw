module MUX13 (MemoryData, SSout, ext16_32, ulaResult, MUX13out)

input [1:0]MemoryData;
input [31:0] SSout, ext16_32, ulaResult, MUX13out;
output [31:0] MUX13out;


