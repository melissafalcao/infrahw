module SighExtend(concatout, ext25_32);

	input muux14; 
	input [25:0]  concatout; 
	output [31:0]  ext25_32;

endmodule
