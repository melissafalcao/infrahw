module SighExtend16_32(imediato, ext16_32);

	input [15:0]  imediato; 
	output [31:0]  ext16_32; 

endmodule
