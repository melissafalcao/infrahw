module MemoryDataRegister(MDR, memoryOut, MDRout) 

input MDR;
input [31:0] memoryOut;
output [31:0] MDRout;