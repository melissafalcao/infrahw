module CONCAT (rs, rt, imediato, concatout);

//concaternar rs,rt e imediato (conferir a ordem da concatenacao, zé n tem certeza)
  input [4:0] rs;
  input [4:0] rt;
  input [15:0] immediato;
output [25:0] concatout;

endmodule
