module LoadSize (LS, MDRout, LSout) 

input [1:0] LS;
input [31:0] MDRout;
output [31:0] LSout;